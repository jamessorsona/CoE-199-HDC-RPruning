parameter integer SHIFTS [0:FEATURE_COUNT-1] = '{
	127,
	536,
	389,
	207,
	72,
	109,
	451,
	124,
	219,
	25,
	520,
	156,
	104,
	349,
	491,
	12,
	181,
	281,
	150,
	437,
	426,
	521,
	473,
	276,
	510,
	293,
	2,
	418,
	407,
	308,
	192,
	602,
	382,
	518,
	543,
	399,
	243,
	502,
	169,
	230,
	591,
	81,
	116,
	336,
	187,
	315,
	33,
	235,
	241,
	292,
	121,
	322,
	376,
	303,
	99,
	277,
	453,
	278,
	412,
	411,
	402,
	32,
	248,
	138,
	261,
	616,
	19,
	445,
	352,
	417,
	202,
	2,
	216,
	483,
	8,
	498,
	375,
	503,
	145,
	265,
	290,
	386,
	80,
	199,
	40,
	507,
	476,
	568,
	46,
	84,
	26,
	479,
	354,
	185,
	454,
	70,
	257,
	489,
	143,
	44,
	268,
	112,
	567,
	419,
	588,
	74,
	182,
	215,
	200,
	226,
	424,
	31,
	173,
	310,
	554,
	43,
	537,
	530,
	516,
	260,
	595,
	500,
	189,
	86,
	488,
	570,
	128,
	279,
	466,
	546,
	519,
	194,
	45,
	436,
	486,
	134,
	95,
	165,
	566,
	288,
	493,
	227,
	211,
	59,
	342,
	413,
	487,
	96,
	56,
	457,
	275,
	250,
	358,
	102,
	328,
	325,
	66,
	272,
	198,
	204,
	434,
	456,
	422,
	448,
	585,
	580,
	409,
	569,
	242,
	381,
	171,
	62,
	37,
	470,
	415,
	323,
	420,
	87,
	14,
	191,
	160,
	430,
	380,
	343,
	151,
	91,
	449,
	129,
	351,
	83,
	224,
	61,
	289,
	439,
	396,
	307,
	529,
	245,
	110,
	259,
	528,
	403,
	228,
	481,
	362,
	298,
	306,
	504,
	427,
	168,
	596,
	478,
	17,
	366,
	1,
	180,
	299,
	218,
	163,
	212,
	16,
	30,
	581,
	397,
	357,
	85,
	111,
	131,
	432,
	93,
	64,
	100,
	274,
	300,
	319,
	459,
	106,
	309,
	592,
	614,
	400,
	355,
	291,
	220,
	206,
	132,
	613,
	540,
	167,
	374,
	373,
	36,
	317,
	541,
	157,
	164,
	152,
	122,
	155,
	238,
	297,
	534,
	222,
	321,
	126,
	414,
	247,
	398,
	367,
	210,
	571,
	232,
	583,
	423,
	597,
	184,
	273,
	589,
	406,
	262,
	7,
	523,
	166,
	610,
	9,
	353,
	431,
	477,
	378,
	316,
	501,
	531,
	421,
	341,
	271,
	78,
	225,
	3,
	379,
	495,
	514,
	320,
	141,
	551,
	98,
	305,
	236,
	393,
	480,
	105,
	564,
	345,
	302,
	371,
	443,
	428,
	555,
	603,
	50,
	544,
	178,
	338,
	162,
	465,
	440,
	186,
	82,
	391,
	363,
	360,
	563,
	365,
	612,
	7,
	217,
	154,
	120,
	287,
	253,
	339,
	532,
	136,
	494,
	333,
	107,
	269,
	574,
	256,
	252,
	474,
	561,
	197,
	71,
	263,
	214,
	130,
	209,
	496,
	246,
	170,
	372,
	312,
	89,
	334,
	284,
	404,
	75,
	575,
	159,
	52,
	505,
	384,
	34,
	125,
	578,
	429,
	395,
	233,
	286,
	295,
	368,
	203,
	401,
	229,
	249,
	55,
	361,
	346,
	579,
	205,
	267,
	76,
	600,
	517,
	49,
	390,
	114,
	142,
	42,
	18,
	285,
	244,
	67,
	188,
	527,
	438,
	133,
	58,
	542,
	25,
	387,
	39,
	329,
	47,
	410,
	140,
	347,
	304,
	364,
	441,
	149,
	559,
	251,
	547,
	506,
	533,
	605,
	221,
	562,
	239,
	35,
	392,
	433,
	594,
	472,
	73,
	196,
	348,
	21,
	565,
	294,
	586,
	377,
	177,
	455,
	388,
	101,
	213,
	599,
	234,
	48,
	223,
	327,
	444,
	350,
	65,
	183,
	356,
	29,
	598,
	485,
	442,
	311,
	65,
	425,
	6,
	201,
	522,
	550,
	4,
	97,
	385,
	557,
	576,
	340,
	463,
	314,
	508,
	53,
	172,
	113,
	359,
	526,
	326,
	509,
	175,
	90,
	601,
	318,
	137,
	266,
	606,
	144,
	68,
	464,
	608,
	615,
	538,
	24,
	313,
	484,
	174,
	416,
	369,
	446,
	176,
	283,
	383,
	103,
	324,
	394,
	147,
	27,
	148,
	41,
	331,
	94,
	604,
	556,
	584,
	408,
	79,
	461,
	558,
	330,
	515,
	54,
	452,
	301,
	190,
	553,
	237,
	549,
	609,
	590,
	255,
	513,
	118,
	545,
	572,
	28,
	462,
	280,
	492,
	270,
	77,
	405,
	135,
	611,
	370,
	607,
	254,
	282,
	115,
	60,
	158,
	1,
	469,
	573,
	161,
	69,
	497,
	475,
	332,
	337,
	460,
	108,
	51,
	490,
	535,
	525,
	435,
	38,
	63,
	117,
	146,
	539,
	88,
	458,
	482,
	153,
	1,
	344,
	587,
	471,
	195,
	512,
	240,
	13,
	524,
	139,
	231,
	123,
	208,
	582,
	467,
	548,
	577,
	593,
	23,
	511,
	560,
	335,
	447,
	552,
	499,
	258,
	17,
	468,
	179,
	1,
	450,
	92,
	264,
	296,
	193,
	119
};
