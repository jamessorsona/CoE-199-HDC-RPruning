`timescale 1ns/1ps
`include "../rtl_wo_rp/am_fsm.sv"
`include "../rtl_wo_rp/am_mux_in.sv"
`include "../rtl_wo_rp/am_and_array.sv"
`include "../rtl_wo_rp/am_tree_adder.sv"
`include "../rtl_wo_rp/am_tree_comparator.sv"
`include "../rtl_wo_rp/class_fsm.sv"
`include "../rtl_wo_rp/class_mux_in.sv"
`include "../rtl_wo_rp/class_bundler.sv"
`include "../rtl_wo_rp/class_thresholder.sv"
`include "../rtl_wo_rp/class_reg_nonbin.sv"
`include "../rtl_wo_rp/class_reg_bin.sv"
`include "../rtl_wo_rp/enc_fsm.sv"
`include "../rtl_wo_rp/enc_binder.sv"
`include "../rtl_wo_rp/enc_nets.sv"
`include "../rtl_wo_rp/enc_mux_in.sv"
`include "../rtl_wo_rp/enc_bundler.sv"
`include "../rtl_wo_rp/enc_reg_out.sv"
`include "../rtl_wo_rp/oneshot_fsm.sv"
`include "../rtl_wo_rp/quantizing_top.sv"
`include "../rtl_wo_rp/encoding_top.sv"
`include "../rtl_wo_rp/class_hv_gen_top.sv"
`include "../rtl_wo_rp/am_top.sv"
`include "../rtl_wo_rp/qtz_fsm.sv"
`include "../rtl_wo_rp/qtz_mux_in.sv"
`include "../rtl_wo_rp/quantizer.sv"
`include "../rtl_wo_rp/qtz_im.sv"
`include "../rtl_wo_rp/qtz_im_fetch.sv"
`include "../rtl_wo_rp/qtz_reg_out.sv"
